// Code your testbench here
// This testbench is tested succesfully on edaplayground

module SR_ff_tb;

reg clk;
reg reset;
reg s,r;

wire q;
wire qb;

sr_ff srflipflop( .clk(clk), .reset(reset), .s(s), .r(r), .q(q), .q_bar(qb) );

initial begin
  $dumpfile("dump.vcd");
  $dumpvars(0,SR_ff_tb);

s = 1'b0;
r = 1'b0;
reset = 1;
clk=1;

#10 
reset=0;
s=1'b1;
r=1'b0;

#100
reset=0;
s=1'b0;
r=1'b1;
#90
  s=1'b0;
  r=1'b0;

#200
  $finish;

end
always #25 clk <= ~clk;

endmodule
